module top(
		output green_led_d7,
		output orange_led_d8,
		output red_led_d5,
		output yellow_led_d6
	);
	assign green_led_d7  = 1;
	assign orange_led_d8 = 1;
	assign red_led_d5    = 1;
	assign yellow_led_d6 = 1;

endmodule
